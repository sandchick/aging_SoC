/*Copyright 2018-2021 T-Head Semiconductor Co., Ltd.

Licensed under the Apache License, Version 2.0 (the "License");
you may not use this file except in compliance with the License.
You may obtain a copy of the License at

    http://www.apache.org/licenses/LICENSE-2.0

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.
*/

module e902_gpio_io();

`define b_pad_porta tb.x_soc.b_pad_gpio_porta[7:0]

initial
begin

  wait(`b_pad_porta == 8'hff);
  $display("************gpio port a output test pass!************");
  
  force `b_pad_porta = 8'hff;
end
endmodule
